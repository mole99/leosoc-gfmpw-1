// SPDX-FileCopyrightText: © 2022 Leo Moser <https://codeberg.org/mole99>
// SPDX-License-Identifier: GPL-3.0-or-later

module arbiter_tb ();
    timeunit 1ns;
    timeprecision 1ps;
endmodule
